module top(
    output      pin
);

assign pin = 1'b1;

endmodule